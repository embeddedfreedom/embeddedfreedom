*Current Mirror with BJT for Early Effect Demo
V1 n1 0 15
RPgm n1 n2 15k
RLoad n1 n3 5k
QPgm n2 n2 0 Q2N3904
QLoad n3 n2 0 Q2N3904

*		Model for 2N3904 NPN BJT (from Eval library in Pspice)
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)

.control
let start_d = 0
let delta_d = 1K
let stop_d = 15K
let d_act = start_d
while d_act le stop_d
     alter RLoad d_act
     echo *****************************
     echo Running sim with RLoad:"$&d_act"
     echo *****************************
     let d_act = d_act + delta_d
     op
     show Qpgm rpgm QLoad rload 
     end
.endc
.end

 